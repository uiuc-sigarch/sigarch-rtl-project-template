//-----------------------------------------------------------------------------
// Title         : SIGARCH Blank Top Test Package
// Project       : SIGARCH Blank RTL
//-----------------------------------------------------------------------------
// File          : sigarch_blank_top_test_pkg.sv
// Author        : Nebhrajani A. V.
// Created       : 21.07.2023
//-----------------------------------------------------------------------------
// Description :
// Top test package for the SIGARCH blank module. Contains all the classes,
// etc. needed by the top level UVM testbench.
//-----------------------------------------------------------------------------
// Copyright (c) SIGARCH@UIUC <sigarch@acm.illinois.edu>
//-----------------------------------------------------------------------------

package sigarch_blank_top_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  // `include "some_agent.svh"
  // ...

endpackage : sigarch_blank_top_test_pkg
